/*
 * Seven-segment display timer for the Minisys board
 */

module mipsfpga_ahb_sevensegtimer(
                     input            clk,
                     input            resetn,
                     input      [7:0] EN,
                     input      [3:0] DISP0,
                     input      [3:0] DISP1,
                     input      [3:0] DISP2,
                     input      [3:0] DISP3,
                     input      [3:0] DISP4,
                     input      [3:0] DISP5,
                     input      [3:0] DISP6,
                     input      [3:0] DISP7,
                     output     [7:0] DISPENOUT,
                     output     [6:0] DISPOUT);

  // Add code here.

endmodule

