/*
 * Seven-segment display decoder
 */

module mipsfpga_ahb_sevensegdec(input      [3:0] data,
                                output reg [6:0] segments);

  // Add code here.

endmodule
